library verilog;
use verilog.vl_types.all;
entity controlAllu_vlg_vec_tst is
end controlAllu_vlg_vec_tst;

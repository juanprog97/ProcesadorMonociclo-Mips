library verilog;
use verilog.vl_types.all;
entity allu_vlg_vec_tst is
end allu_vlg_vec_tst;

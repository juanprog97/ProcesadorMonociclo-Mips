library verilog;
use verilog.vl_types.all;
entity registrosFicheros_vlg_vec_tst is
end registrosFicheros_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity programCounter_vlg_vec_tst is
end programCounter_vlg_vec_tst;

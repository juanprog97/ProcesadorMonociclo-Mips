library verilog;
use verilog.vl_types.all;
entity unidadControl_vlg_vec_tst is
end unidadControl_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity MIPS is
    port(
        Clock           : in     vl_logic
    );
end MIPS;

library verilog;
use verilog.vl_types.all;
entity memoriaRam_vlg_vec_tst is
end memoriaRam_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity multiplexor_vlg_vec_tst is
end multiplexor_vlg_vec_tst;

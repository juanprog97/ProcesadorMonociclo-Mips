library verilog;
use verilog.vl_types.all;
entity memoriaInstrucciones_vlg_vec_tst is
end memoriaInstrucciones_vlg_vec_tst;
